module directory

pub enum SearchOption {
	top_only
	recursive
}
